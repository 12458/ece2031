-- IO DECODER for SCOMP
-- This eliminates the need for a lot of AND decoders or Comparators 
--    that would otherwise be spread around the top-level BDF

LIBRARY IEEE;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY IO_DECODER IS
  PORT (
    IO_ADDR       : IN  STD_LOGIC_VECTOR(10 downto 0);
    IO_CYCLE      : IN  STD_LOGIC;

    SWITCH_EN     : OUT STD_LOGIC;
    TIMER_EN      : OUT STD_LOGIC;
    HEX0_EN       : OUT STD_LOGIC;
    HEX1_EN       : OUT STD_LOGIC;

    LED_TOGGLE_EN     : OUT STD_LOGIC;
    LED_BRIGHTNESS_EN : OUT STD_LOGIC;
    LED_EFFECTS_EN    : OUT STD_LOGIC;

    LED_INDEX_VECTOR  : OUT STD_LOGIC_VECTOR(9 downto 0)
  );
END ENTITY;


ARCHITECTURE a OF IO_DECODER IS
  SIGNAL ADDR_INT : INTEGER RANGE 0 TO 2047;
BEGIN

  ADDR_INT <= TO_INTEGER(UNSIGNED(IO_ADDR));

  SWITCH_EN <= '1' WHEN (ADDR_INT = 16#000#) AND (IO_CYCLE = '1') ELSE '0';
  TIMER_EN  <= '1' WHEN (ADDR_INT = 16#002#) AND (IO_CYCLE = '1') ELSE '0';
  HEX0_EN   <= '1' WHEN (ADDR_INT = 16#004#) AND (IO_CYCLE = '1') ELSE '0';
  HEX1_EN   <= '1' WHEN (ADDR_INT = 16#005#) AND (IO_CYCLE = '1') ELSE '0';

  LED_TOGGLE_EN     <= '1' WHEN (ADDR_INT = 16#020#) AND (IO_CYCLE = '1') ELSE '0';
  LED_BRIGHTNESS_EN <= '1' WHEN (ADDR_INT = 16#021#) AND (IO_CYCLE = '1') ELSE '0';
  LED_EFFECTS_EN    <= '1' WHEN (ADDR_INT = 16#02C#) AND (IO_CYCLE = '1') ELSE '0';

  LED_INDEX_VECTOR <= 
    "0000000001" WHEN (ADDR_INT = 16#022#) AND (IO_CYCLE = '1') ELSE
    "0000000010" WHEN (ADDR_INT = 16#023#) AND (IO_CYCLE = '1') ELSE
    "0000000100" WHEN (ADDR_INT = 16#024#) AND (IO_CYCLE = '1') ELSE
    "0000001000" WHEN (ADDR_INT = 16#025#) AND (IO_CYCLE = '1') ELSE
    "0000010000" WHEN (ADDR_INT = 16#026#) AND (IO_CYCLE = '1') ELSE
    "0000100000" WHEN (ADDR_INT = 16#027#) AND (IO_CYCLE = '1') ELSE
    "0001000000" WHEN (ADDR_INT = 16#028#) AND (IO_CYCLE = '1') ELSE
    "0010000000" WHEN (ADDR_INT = 16#029#) AND (IO_CYCLE = '1') ELSE
    "0100000000" WHEN (ADDR_INT = 16#02A#) AND (IO_CYCLE = '1') ELSE
    "1000000000" WHEN (ADDR_INT = 16#02B#) AND (IO_CYCLE = '1') ELSE
    (others => '0');

END a;
